
module hazard_detection_unit (
    input logic i_clk,
    input logic i_reset,
    
    // Register dependencies
    input logic [4:0] i_id_rs1,          // Source register 1 in ID stage
    input logic [4:0] i_id_rs2,          // Source register 2 in ID stage
    input logic [4:0] i_ex_rd,           // Destination register in EX stage
    input logic [4:0] i_mem_rd,          // Destination register in MEM stage
    
    // Instruction types
    input logic i_ex_mem_read,            // Load instruction in EX stage
    // input logic i_ex_reg_write,           // Register write in EX stage
    // input logic i_mem_reg_write,          // Register write in MEM stage
    
    // Branch/jump detection
    input logic i_branch_taken,           // Branch taken signal
    input logic i_jump_taken,             // Jump taken signal
    
    // Hazard outputs
    output logic o_stall,                 // Stall pipeline
    output logic o_flush                  // Flush pipeline stages
);

    // 1. Load-use data hazards
    // 2. Control hazards (branches/jumps)
    // 3. Structural hazards
    
    always_comb begin
        o_stall = 1'b0;
        o_flush = 1'b0;

        // control hazards 
        if (i_branch_taken || i_jump_taken) begin
            o_flush = 1'b1;
        end
        
        // load-use hazards
        else if (i_ex_mem_read && 
            ((i_ex_rd == i_id_rs1) || (i_ex_rd == i_id_rs2)) &&
            (i_ex_rd != 5'b0)) begin
            o_stall = 1'b1;
        end
    end

endmodule
