module alu_control (
    
);
    
endmodule
