`ifndef CONFIG_H
`define CONFIG_H

`define USE_ROM
// `define USE_STATIC
`define SHOW_INITIAL_MEMORY

`define PROGRAM_FILE "mem/test_rv32i.hex"

`endif //CONFIG_H
