`define WIDTH 32

module top (
    input logic clk,
    input logic reset 
);
    
endmodule
