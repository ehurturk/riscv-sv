`define ALU_OPSIZE 4
