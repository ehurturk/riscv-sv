// Pipelined datapath

module pipelined_datapath (
    input logic clk,
    input logic reset
);



endmodule
