`ifndef CONFIG_H
`define CONFIG_H

`define USE_ROM
// `define USE_STATIC
`define SHOW_INITIAL_MEMORY

`define PROGRAM_FILE "mem/test_simple_br.hex"
// `define PROGRAM_FILE "mem/test_br.hex"

`endif //CONFIG_H
