// multi cycle control unit FSM


module mccontrol (
    
);
    
endmodule : mccontrol
