module regfile (
    ports 
    input logic write_enable;
    output logic [31:0] r_data1;
    output logic [31:0] r_data2;
);
    
endmodule