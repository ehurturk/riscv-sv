`ifndef CONFIG_H
`define CONFIG_H

`define USE_ROM
// `define USE_STATIC
`define SHOW_INITIAL_MEMORY

`endif //CONFIG_H
